module day5(input x, input y, output z);
  xnor(z,x,y);
endmodule
